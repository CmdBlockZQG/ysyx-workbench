typedef enum {
  PERF_IFU_FETCH,
  PERF_IDU_UPIMM,
  PERF_IDU_JUMP,
  PERF_IDU_BRANCH,
  PERF_IDU_LOAD,
  PERF_IDU_STORE,
  PERF_IDU_CALRI,
  PERF_IDU_CALRR,
  PERF_IDU_SYS,
  PERF_IDU_CSR,
  PERF_EXU_UPIMM,
  PERF_EXU_JUMP,
  PERF_EXU_BRANCH,
  PERF_EXU_LOAD,
  PERF_EXU_STORE,
  PERF_EXU_CALRI,
  PERF_EXU_CALRR,
  PERF_EXU_SYS,
  PERF_EXU_CSR,
  PERF_EXU_READY,
  PERF_LSU_LOAD,
  PERF_LSU_LOAD_RESP,
  PERF_LSU_WRITE
} perf_cnt_t;
