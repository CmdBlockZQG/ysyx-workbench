// 访存Funct常量
parameter reg [2:0] LD_BS = 3'b000;
parameter reg [2:0] LD_HS = 3'b001;
parameter reg [2:0] LD_W  = 3'b010;
parameter reg [2:0] LD_BU = 3'b100;
parameter reg [2:0] LD_HU = 3'b101;

parameter reg [2:0] ST_B = 3'b000;
parameter reg [2:0] ST_H = 3'b001;
parameter reg [2:0] ST_W = 3'b010;
