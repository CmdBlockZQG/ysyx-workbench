typedef enum {
  PERF_IFU_FETCH,
  PERF_LSU_LOAD_RESP,
  PERF_EXU_READY,
  PERF_IDU_UPIMM,
  PERF_IDU_JUMP,
  PERF_IDU_BRANCH,
  PERF_IDU_LOAD,
  PERF_IDU_STORE,
  PERF_IDU_CALRI,
  PERF_IDU_CALRR,
  PERF_IDU_SYS,
  PERF_IDU_CSR
} perf_cnt_t;
