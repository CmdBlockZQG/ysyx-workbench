// Branch指令Funct常量
parameter BR_BEQ  = 3'b000;
parameter BR_BNE  = 3'b001;
parameter BR_BLT  = 3'b100;
parameter BR_BGE  = 3'b101;
parameter BR_BLTU = 3'b110;
parameter BR_BGEU = 3'b111;
