typedef enum {
  PERF_IFU_WAIT,
  PERF_IFU_INST,
  PERF_IFU_HOLD,
  PERF_ICACHE_MISS,
  PERF_ICACHE_MEM,
  PERF_IDU_IDLE,
  PERF_IDU_INST,
  PERF_IDU_HOLD,
  PERF_IDU_LOAD,
  PERF_IDU_STORE,
  PERF_IDU_BRANCH,
  PERF_IDU_JAL,
  PERF_IDU_JALR,
  PERF_EXU_IDLE,
  PERF_EXU_INST,
  PERF_EXU_FLUSH,
  PERF_EXU_MEMR,
  PERF_EXU_MEMW
} perf_cnt_t;
