// 访存Funct常量
parameter LD_BS = 3'b000;
parameter LD_HS = 3'b001;
parameter LD_W  = 3'b010;
parameter LD_BU = 3'b100;
parameter LD_HU = 3'b101;

parameter ST_B = 3'b000;
parameter ST_H = 3'b001;
parameter ST_W = 3'b010;
