typedef enum {
  PERF_IFU_FETCH,
  PERF_IFU_WAIT_MEM,
  PERF_IFU_WAIT_EXU,
  PERF_IDU_UPIMM,
  PERF_IDU_JUMP,
  PERF_IDU_BRANCH,
  PERF_IDU_LOAD,
  PERF_IDU_STORE,
  PERF_IDU_CALRI,
  PERF_IDU_CALRR,
  PERF_IDU_SYS,
  PERF_IDU_CSR,
  PERF_EXU_UPIMM,
  PERF_EXU_JUMP,
  PERF_EXU_BRANCH,
  PERF_EXU_LOAD,
  PERF_EXU_STORE,
  PERF_EXU_CALRI,
  PERF_EXU_CALRR,
  PERF_EXU_SYS,
  PERF_EXU_CSR,
  PERF_EXU_READY,
  PERF_LSU_LOAD,
  PERF_LSU_LOAD_RESP,
  PERF_LSU_STORE,
  PERF_ICACHE_HIT,
  PERF_ICACHE_MISS,
  PERF_ICACHE_WAIT_MEM
} perf_cnt_t;
