// opcode 常量
parameter OP_LUI    = 5'b01101;
parameter OP_AUIPC  = 5'b00101;
parameter OP_JAL    = 5'b11011;
parameter OP_JALR   = 5'b11001;
parameter OP_BRANCH = 5'b11000;
parameter OP_LOAD   = 5'b00000;
parameter OP_STORE  = 5'b01000;
parameter OP_CALRI  = 5'b00100;
parameter OP_CALRR  = 5'b01100;
parameter OP_SYS    = 5'b11100;
